module test(input clk);
    logic[12:0] v,w;
    // assign v[3:0] = 32'b0;
    // assign w[4:0] = 32'b0;
endmodule