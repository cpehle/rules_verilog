module test_2(input clk);
    logic[12:0] v;
    // assign v[3:0] = 32'b0;
endmodule